//module NNAccelerator